// no timescale needed

module conv_std_logic_vector_demo(
input wire [7:0] x,
output wire [7:0] y
);





  // triggers two-argument conv_std_logic_vector usage
  assign y = (5) ^ x;

endmodule
