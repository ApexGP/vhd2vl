// no timescale needed

module concat_demo(
input wire reset
);

parameter [26:0] abc={3'b010,12'haaa};
parameter [31:0] xyz=32'h000000ff;




endmodule  // incomplete: entity-only
